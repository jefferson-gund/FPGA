-- Rom de imagem do objeto "POU"

library ieee;
use ieee.std_logic_1164.all;
library work;
use work.vga_package.all;

entity pou_rom is
	
	port
	(
		-- Input ports
		x_pou : in integer range 0 to hpou;
		y_pou : in integer range 0 to vpou;

		-- Output ports
		rgb_pou : out std_logic_vector(2 downto 0)
	);
end pou_rom;

architecture estrutura of pou_rom is
	
	constant POU : matrix_pou :=(
			
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","011","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","111","111","111","011","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","011","011","011","011","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","001","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","011","011","111","111","111","111","111","111","111","111","111","111","111","011","011","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","011","011","011","011","011","001","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","011","011","011","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","011","011","000","011","011","011","011","011","011","011","011","011","011","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","011","011","011","011","011","011","011","011","011","001","001","011","011","001","001","001","001","001","000","000","000","000","000","001","001","001","001","000","001","111","111","111","111","111","111","111","111","111","111","001","011","011","011","011","011","011","011","011","011","011","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","001","011","011","011","011","011","011","011","011","011","001","111","111","111","111","111","111","111","111","111","111","111","111","001","011","011","011","011","011","111","111","111","111","111","111","111","111","111","111","111","111","001","011","011","011","011","011","011","011","011","011","001","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","011","011","011","011","011","011","011","011","011","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","011","011","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","011","011","011","011","011","011","011","011","011","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","011","011","011","011","011","011","011","011","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","011","011","011","011","011","011","011","011","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","011","011","011","011","011","011","011","011","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","011","011","011","011","011","011","011","011","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","011","011","011","011","011","011","011","011","001","111","111","111","111","111","111","001","000","000","001","111","111","111","111","111","111","001","001","111","111","111","111","111","111","001","000","000","001","111","111","111","111","111","111","001","011","011","011","011","011","011","011","011","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","011","011","011","011","011","011","011","011","011","111","111","111","111","111","001","000","000","000","000","001","111","111","111","111","111","001","011","111","111","111","111","111","001","000","000","000","000","001","111","111","111","111","111","011","011","011","011","011","011","011","011","011","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","011","001","000","000","000","011","011","011","011","011","011","011","011","011","111","111","111","111","111","000","000","000","000","000","000","111","111","111","111","111","011","011","111","111","111","111","111","000","000","000","000","000","000","111","111","111","111","111","011","011","011","011","011","011","011","011","011","000","000","000","001","011","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","011","011","001","000","000","000","011","011","011","011","011","011","011","011","011","111","111","111","111","111","001","000","000","000","000","001","111","111","111","111","111","001","011","111","111","111","111","111","001","000","000","000","000","001","111","111","111","111","111","011","011","011","011","011","011","011","011","011","000","000","000","001","011","011","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","011","011","011","000","000","000","001","011","011","011","011","011","011","011","001","111","111","111","111","111","111","001","000","000","000","111","111","111","111","111","111","001","001","111","111","111","111","111","111","000","000","000","001","111","111","111","111","111","111","001","011","011","011","011","011","011","011","001","000","000","000","011","011","011","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","011","011","011","011","000","000","000","001","011","011","011","011","011","011","011","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","011","011","011","011","011","011","011","001","000","000","000","011","011","011","011","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","011","011","011","011","011","001","000","000","000","011","011","011","011","011","011","011","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","011","011","011","011","011","011","011","000","000","000","001","011","011","011","011","011","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","001","000","000","000","011","011","011","011","011","011","011","011","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","011","011","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","011","011","011","011","011","011","011","011","000","000","000","001","011","011","011","011","011","011","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","011","000","000","000","000","011","011","011","011","011","011","011","001","001","111","111","111","111","111","111","111","111","111","111","111","111","011","001","000","000","001","011","111","111","111","111","111","111","111","111","111","111","111","111","011","011","011","011","011","011","011","011","011","000","000","000","000","011","011","011","011","011","011","011","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","001","000","000","000","001","011","011","011","011","011","011","011","001","011","111","111","111","111","111","111","111","111","111","111","011","001","001","000","000","001","001","011","111","111","111","111","111","111","111","111","111","111","011","001","011","011","011","011","011","011","011","001","000","000","000","001","011","011","011","011","011","011","011","011","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","000","000","000","000","001","011","011","011","011","011","011","011","011","001","111","111","111","111","111","111","111","111","001","001","001","000","000","000","000","001","001","001","111","111","111","111","111","111","111","111","001","011","011","011","011","011","011","011","011","001","000","000","000","000","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","000","000","000","000","000","001","011","011","011","011","011","011","011","011","001","001","001","001","001","001","001","001","000","000","000","001","001","000","000","000","001","001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","001","000","000","000","000","000","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","001","000","000","000","000","000","000","001","001","001","011","011","011","011","011","001","001","000","000","000","000","000","000","011","011","011","011","000","000","000","000","000","000","001","001","011","011","011","011","011","001","001","001","000","000","000","000","000","000","001","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","011","011","011","011","011","011","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","000","000","000","000","000","000","000","000","000","000","000","000","001","011","011","011","011","011","011","011","011","011","011","011","011","001","000","000","000","000","000","000","000","000","000","000","000","000","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001","001"),
			("001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001","001"),
			("001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001"),
			("001","001","001","001","001","111","111","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","111","111","111","001","001","001","001","001"),
			("001","001","001","001","111","111","111","111","111","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","111","111","111","111","111","111","001","001","001","001"),
			("001","001","001","001","111","111","111","111","111","111","111","111","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","000","000","000","000","000","000","000","000","000","000","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","111","111","111","111","111","111","111","111","001","001","001","001"),
			("001","001","001","000","001","111","111","111","111","111","111","111","111","111","111","111","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","000","000","000","000","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","111","111","111","111","111","111","111","111","111","111","111","000","000","001","001","001"),
			("001","001","001","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","111","111","111","111","111","111","111","111","111","111","111","111","111","001","000","000","000","001","001","001"),
			("001","001","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","000","000","000","000","000","000","001","001"),
			("001","001","000","000","000","000","000","000","000","000","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","011","011","011","011","011","011","011","011","011","011","001","001","011","011","011","011","011","011","011","011","011","001","001","001","011","011","011","011","011","011","011","011","011","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","000","000","000","000","000","000","000","000","001","001"),
			("001","000","000","000","000","000","000","000","000","000","000","000","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001","011","011","011","011","001","001","001","001","001","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","000","000","000","000","000","000","000","000","000","000","000","000","001"),
			("001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001"),
			("001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001"),
			("001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001"),
			("001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","011","011","011","111","111","111","111","111","111","001","001","001","001","001","111","111","001","111","111","111","001","001","001","001","101","111","111","111","111","111","111","011","011","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001"),
			("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","111","111","001","001","111","111","111","111","111","111","111","111","111","101","001","001","111","111","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000"),
			("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","111","111","111","111","111","111","111","111","111","111","111","111","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000"),
			("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","111","111","111","111","111","111","111","111","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000"),
			("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000"),
			("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000"),
			("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000"),
			("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000"),
			("000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000"),
			("001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001"),
			("001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","101","101","101","101","101","101","101","101","101","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001"),
			("001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001"),
			("001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","111","111","111","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001"),
			("001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001"),
			("001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001"),
			("001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001"),
			("001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001"),
			("001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","111","111","111","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001"),
			("001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","111","111","111","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","111","111","111","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","011","111","011","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001")
	);
											
begin

	rgb_pou <= POU(y_pou,x_pou);

end estrutura;
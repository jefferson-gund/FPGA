library ieee;
use ieee.std_logic_1164.all;
library work;
use work.vga_package.all;

entity play_symbols is
	
	port
	(
		-- Input ports
		index : in integer range 0 to 2;
		x_play : in integer range 0 to hplay;
		y_play : in integer range 0 to vplay;
		-- Output ports
		rgb_colour : out std_logic_vector(2 downto 0) 

	);
end play_symbols;

architecture lista of play_symbols is
	
	constant start : matrix_play :=(
			
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001","001","001","001","001"),
			("001","001","001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001","001","001"),
			("001","001","001","001","001","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001","001","001"),
			("001","001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","011","001","001","001"),
			("001","001","001","001","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001","001"),
			("001","001","001","011","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","110","100","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","110","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","110","100","110","110","110","110","100","100","100","100","100","100","100","110","110","110","100","110","110","100","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","110","100","100","100","110","110","110","100","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","110","110","100","100","100","100","110","110","110","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","100","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","100","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","100","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","110","110","110","110","110","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","100","100","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","100","100","100","100","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","100","100","100","100","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","100","100","100","100","110","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","100","100","100","100","110","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","100","100","100","100","100","100","100","100","100","100","110","110","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","001","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001","001"),
			("001","001","001","001","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001","001"),
			("001","001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001","001"),
			("001","001","001","001","001","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001","001","001"),
			("001","001","001","001","001","011","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001","001","001","001"),
			("001","001","001","001","001","001","011","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001")
	);

















		constant pause : matrix_play :=(
		
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","001","001","001","001","001","001"),
			("001","001","001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001","001","001"),
			("001","001","001","001","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","110","110","110","110","110","110","110","100","100","100","100","100","100","100","110","110","110","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","100","100","100","100","100","110","100","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","100","100","100","100","100","110","100","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","100","100","100","100","100","110","100","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","100","100","100","100","100","110","100","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","110","110","110","110","110","110","110","100","110","110","110","110","110","110","110","110","110","110","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","110","100","110","110","100","100","100","100","100","100","110","110","110","110","100","100","100","110","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","110","110","110","110","110","110","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","100","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","100","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","110","100","110","110","110","110","110","110","110","110","100","100","100","100","100","100","100","100","100","100","100","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001"),
			("001","001","011","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001"),
			("001","001","001","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001"),
			("001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","001","001","001"),
			("001","001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","011","001","001","001"),
			("001","001","001","001","001","111","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","110","111","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001")
	);






	
	constant game_over : matrix_play :=(
	
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001"),
			("001","001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001"),
			("001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001"),
			("001","001","001","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001"),
			("001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001"),
			("001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","111","101","100","100","111","111","111","111","111","111","111","111","111","111","101","100","100","111","111","111","111","111","111","111","111","111","111","111","101","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","101","111","111","111","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","101","111","111","111","111","101","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","100","100","100","100","100","100","100","100","100","100","101","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","101","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","101","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","111","111","111","111","101","100","100","100","111","111","111","111","111","111","111","111","111","111","111","101","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","101","100","101","101","101","100","101","101","101","101","101","101","101","101","111","111","111","111","111","111","111","111","111","111","101","101","101","101","111","111","111","111","111","111","111","111","111","101","101","100","101","111","111","111","111","111","111","111","111","111","111","101","101","101","111","111","111","101","101","101","100","101","101","101","101","101","101","101","101","111","111","111","111","111","111","111","111","100","101","101","101","101","101","101","101","101","101","101","101","101","111","111","111","111","111","100","100","101","111","111","111","111","111","111","111","111","111","101","101","101","101","111","111","111","101","101","101","101","101","101","101","101","101","101","101","101","111","111","101","101","101","101","101","101","101","101","101","101","101","101","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","101","100","100","100","100","111","111","111","111","111","111","111","111","111","100","100","100","100","111","111","111","111","111","111","111","111","111","100","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","101","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","100","100","100","100","100","100","100","100","100","100","100","100","101","111","111","001"),
			("001","001","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","100","100","100","100","100","111","111","111","111","111","111","111","111","111","100","100","100","100","111","111","111","111","111","111","111","111","111","100","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","101","100","100","100","100","100","100","100","100","100","100","100","100","100","100","101","111","111","101","100","100","100","111","111","111","111","111","111","111","111","111","100","100","100","101","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","100","100","100","100","100","100","100","100","100","100","100","100","101","111","111","001"),
			("001","001","111","111","111","111","101","101","101","101","101","101","101","101","101","101","101","101","101","101","111","111","111","111","111","111","111","111","111","111","101","101","111","101","111","111","111","111","111","111","111","111","111","111","101","101","101","111","111","111","111","111","111","111","111","111","101","111","111","101","111","111","111","101","101","100","101","101","101","101","101","101","101","101","101","111","111","111","111","111","111","111","111","101","101","101","101","101","101","101","101","101","101","101","111","101","101","111","111","111","111","101","101","111","111","111","111","111","111","111","111","111","111","101","101","111","111","111","111","111","101","101","100","101","101","101","101","101","101","101","101","101","111","111","101","101","101","101","101","101","101","101","101","101","111","101","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","101","101","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","100","101","101","100","111","111","111","111","111","111","111","111","111","101","100","100","100","101","111","111","111","111","111","111","111","111","101","101","101","101","111","111","111","101","100","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","111","111","111","111","101","101","101","111","111","111","101","101","100","101","111","111","111","111","111","111","111","111","100","101","101","111","111","111","111","101","100","100","111","111","111","111","111","111","111","111","111","111","111","101","100","100","111","111","111","111","111","111","111","101","100","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","100","100","100","111","111","111","111","111","111","111","111","111","101","100","100","100","100","111","111","111","111","111","111","111","111","100","100","100","100","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","100","100","100","100","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","101","100","100","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","100","100","100","100","100","111","111","111","111","111","111","111","111","100","100","100","100","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","100","100","100","100","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","101","100","100","111","111","111","001"),
			("001","001","111","111","111","111","101","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","101","101","101","101","111","111","111","111","111","111","111","111","111","101","100","101","101","101","111","111","111","111","111","111","111","111","101","101","101","101","111","111","111","101","100","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","111","111","111","111","101","101","101","111","111","111","101","100","101","101","111","111","111","111","111","111","111","111","101","101","101","111","111","111","111","101","100","101","111","111","111","111","111","111","111","111","111","111","111","101","100","101","111","111","111","111","111","111","111","101","101","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","101","101","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","101","101","111","101","101","101","101","111","111","111","111","111","111","111","101","101","101","101","101","111","111","111","111","111","111","111","101","101","101","101","101","111","111","111","101","101","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","101","111","111","111","111","111","111","111","111","111","111","101","101","101","111","111","111","111","101","101","101","111","111","111","111","111","111","111","101","101","111","111","111","111","111","111","101","101","101","111","111","111","111","111","111","111","111","111","111","111","101","101","101","111","111","111","111","111","111","111","100","101","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","100","101","100","100","100","100","111","111","111","111","111","111","111","100","100","100","100","100","101","111","111","111","111","111","101","100","100","100","100","100","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","100","100","100","101","111","111","111","111","111","101","100","100","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","101","100","100","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","100","111","101","100","100","100","111","111","111","111","111","111","111","100","100","100","100","100","100","111","111","111","111","111","101","100","100","100","100","100","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","100","100","100","100","111","111","111","111","111","101","100","100","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","101","100","100","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","100","111","111","100","100","101","111","111","111","111","111","111","111","100","100","100","100","100","100","111","111","111","111","111","101","100","100","101","101","100","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","101","100","100","101","111","111","111","111","111","101","100","100","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","101","100","100","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","101","100","100","111","111","111","101","100","100","100","100","100","100","100","101","111","111","111","111","111","111","100","100","101","111","111","111","101","101","101","111","111","111","111","111","111","111","101","100","100","100","100","100","111","111","111","111","111","101","101","101","101","101","101","111","111","111","100","100","100","100","100","100","100","101","101","101","100","101","111","111","111","111","111","111","111","111","100","100","111","111","111","111","111","111","111","111","111","111","101","101","101","111","111","111","111","111","100","100","100","111","111","111","111","111","101","101","100","111","111","111","111","111","111","101","100","100","100","100","100","100","101","101","101","100","101","111","111","101","100","100","101","100","100","100","100","100","100","101","100","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","101","100","100","100","100","100","100","100","100","111","111","111","111","111","111","100","100","100","111","111","111","100","100","100","101","111","111","111","111","111","111","100","100","100","100","100","100","101","111","111","111","111","100","100","100","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","100","100","100","101","111","111","111","101","100","100","100","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","101","100","100","100","100","100","100","100","100","111","111","111","111","111","101","100","100","100","111","111","111","100","100","100","100","111","111","111","111","111","111","100","100","100","100","100","100","101","111","111","111","111","100","100","100","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","100","100","100","101","111","111","111","101","100","100","100","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","101","100","100","100","100","100","100","100","100","111","111","111","111","111","101","100","100","101","111","111","111","101","100","100","100","111","111","111","111","111","111","100","100","100","100","100","100","111","111","111","111","101","100","100","100","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","101","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","100","100","100","101","111","111","111","101","100","100","100","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","001"),
			("001","001","111","111","111","111","101","101","101","111","111","111","111","101","111","111","111","111","111","101","111","111","111","111","111","111","111","101","101","111","111","111","111","111","101","101","101","111","111","111","111","111","111","111","101","101","101","100","100","111","111","111","111","111","101","111","111","111","101","101","111","111","111","100","101","101","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","101","101","111","111","111","111","101","101","101","111","111","111","111","111","111","111","100","100","101","101","111","101","111","111","111","111","111","111","111","111","101","101","101","101","101","101","101","101","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","101","100","101","111","111","111","111","111","111","111","111","111","111","101","101","111","111","111","111","111","101","101","101","111","111","111","111","111","111","101","101","111","111","111","111","111","111","101","101","101","101","100","100","100","111","111","111","100","100","111","111","101","101","101","111","111","111","100","100","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","111","111","111","111","111","111","111","111","111","111","101","101","101","111","111","111","111","111","111","101","101","101","111","111","111","100","101","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","111","111","111","111","111","111","100","101","101","111","101","100","101","101","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","100","100","111","111","111","111","111","100","100","100","101","111","111","111","111","101","100","100","111","111","111","111","111","111","100","100","100","100","100","100","100","101","111","111","100","100","101","111","101","100","100","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","101","100","100","100","111","111","111","100","100","101","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","101","100","100","100","100","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","100","100","111","111","111","111","101","100","100","100","101","111","111","111","111","101","100","100","111","111","111","111","111","111","100","100","100","101","100","100","100","101","111","101","100","100","101","111","101","100","100","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","111","100","100","100","101","111","111","100","100","101","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","100","100","100","100","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","100","100","111","111","111","111","101","100","100","100","111","111","111","111","111","101","100","100","111","111","111","111","111","111","100","100","100","101","100","100","100","101","111","101","100","100","101","111","101","100","100","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","111","100","100","100","101","111","111","100","100","101","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","101","100","100","100","101","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","101","100","100","111","111","111","111","111","111","111","111","111","111","100","101","111","111","111","111","101","100","100","101","111","111","111","111","111","101","101","101","111","111","111","111","111","111","101","100","100","111","101","100","100","101","111","111","100","100","111","111","101","100","101","111","111","111","100","100","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","111","111","111","111","111","111","111","111","111","111","101","101","101","111","111","111","111","111","111","100","100","100","101","111","111","100","100","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","100","100","100","101","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","100","100","111","111","111","111","100","100","100","111","101","100","101","101","100","101","100","100","101","111","111","111","111","111","100","100","100","111","111","100","100","101","111","101","100","100","111","111","101","100","100","111","111","111","100","100","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","111","111","111","111","100","101","101","111","111","111","111","111","111","101","100","100","100","111","101","100","100","101","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","101","100","100","100","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","100","100","111","111","111","111","100","100","100","101","100","100","100","100","100","100","100","100","100","101","111","111","111","111","100","100","100","111","111","100","100","100","111","100","100","100","111","111","101","100","100","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","111","101","100","100","100","100","100","100","100","101","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","101","100","100","100","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","100","100","111","111","111","101","100","100","100","100","100","100","100","100","100","100","100","100","100","101","111","111","111","111","100","100","100","111","111","100","100","100","101","100","100","100","111","111","101","100","100","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","111","111","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","100","100","100","101","111","111","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","100","100","111","111","111","101","100","100","100","100","100","100","100","100","100","100","100","100","100","101","111","111","111","111","100","100","100","111","111","100","100","100","101","100","100","100","111","111","101","100","100","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","111","111","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","100","100","100","100","111","111","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","100","100","111","111","111","101","100","100","100","101","100","100","100","101","101","100","101","100","100","101","111","111","111","111","100","100","100","111","111","100","100","100","101","100","100","101","111","111","101","100","100","111","111","111","100","100","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","111","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","111","111","100","100","100","100","100","100","101","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","101","100","100","100","111","111","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","101","100","100","111","111","111","100","100","100","101","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","100","100","100","111","111","101","100","100","100","100","100","111","111","111","101","100","100","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","111","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","111","111","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","100","100","100","101","111","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","100","100","100","101","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","100","100","100","111","111","101","100","100","100","100","100","111","111","111","100","100","100","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","100","100","100","101","111","111","111","111","111","111","111","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","100","100","100","101","111","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","101","111","111","111","111","111","111","111","101","100","100","100","111","111","101","100","100","100","101","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","100","100","100","111","111","101","100","100","100","100","100","111","111","111","101","100","100","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","100","100","100","101","111","111","111","111","111","111","111","101","100","100","100","100","100","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","111","100","100","100","100","111","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","101","100","100","100","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","100","100","100","111","111","111","100","100","100","100","100","111","111","111","101","100","100","111","111","101","100","100","100","100","100","100","100","100","100","100","100","101","111","111","111","111","111","111","111","101","100","100","100","100","100","100","100","100","100","100","100","100","100","100","101","111","111","111","111","111","111","111","101","100","100","100","100","100","111","111","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","101","111","111","100","100","100","111","111","111","111","111","100","100","100","101","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","101","100","100","100","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","100","100","100","111","111","111","101","100","100","100","100","111","111","111","101","100","101","111","111","111","100","100","100","100","100","100","100","100","100","100","100","101","111","111","111","111","111","111","111","101","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","100","100","100","100","100","111","111","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","101","111","111","100","100","100","111","111","111","111","111","100","100","100","100","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","101","100","100","101","111","111","111","111","111","111","111","111","111","100","100","100","101","111","111","111","100","100","100","111","111","111","101","100","100","100","101","111","111","111","101","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","101","111","111","111","111","111","111","111","101","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","111","101","100","100","100","101","111","111","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","100","100","100","111","111","111","111","111","100","100","100","100","111","111","111","001"),
			("001","001","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","100","100","100","101","111","111","111","111","111","111","111","111","111","100","100","100","100","111","111","111","100","100","100","111","111","111","101","100","100","100","101","111","111","111","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","101","111","111","111","111","111","111","111","101","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","111","101","100","100","100","101","111","111","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","100","100","100","111","111","111","111","111","101","100","100","100","111","111","111","001"),
			("001","001","111","111","111","111","101","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","100","100","100","101","111","111","111","111","111","111","111","111","111","101","100","100","100","111","111","111","100","100","100","111","111","111","101","100","100","100","101","111","111","111","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","101","111","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","111","101","100","100","100","101","111","111","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","100","100","100","111","111","111","111","111","111","100","100","100","101","111","111","001"),
			("001","001","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","101","111","111","101","100","100","100","101","111","111","111","111","111","111","111","111","111","111","100","100","100","111","111","111","100","100","100","111","111","111","101","100","100","100","111","111","111","111","100","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","101","111","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","111","101","100","100","100","111","111","111","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","111","111","100","100","100","111","111","111","111","111","111","100","100","100","100","111","111","001"),
			("001","001","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","100","101","111","111","101","100","100","100","111","111","111","111","111","111","111","111","111","111","111","101","100","100","111","111","111","100","100","100","111","111","111","111","100","100","100","111","111","111","111","101","100","100","111","111","111","100","100","100","100","100","100","100","100","100","100","100","101","111","111","111","111","111","111","111","111","101","100","100","100","100","100","100","100","100","100","100","100","100","111","111","111","111","111","111","111","111","111","111","111","100","100","101","111","111","111","111","111","111","111","111","111","111","100","100","100","100","100","100","100","100","100","100","100","101","111","111","100","100","100","111","111","111","111","111","111","101","100","100","100","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","101","111","111","111","101","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","101","101","111","111","111","111","111","111","111","111","101","101","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001"),
			("001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","001"),
			("001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001"),
			("001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001"),
			("001","001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001"),
			("001","001","001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001")
	);

















											
begin

	rgb_colour <= start(y_play,x_play) 				when index = 0 else
					  pause(y_play,x_play) 				when index = 1 else
					  game_over(y_play,x_play) 		when index = 2 else
					  "000";
end lista;
-- Rom de Figuras Padrão 30 x 30

library ieee;
use ieee.std_logic_1164.all;
library work;
use work.vga_package.all;

entity rom_symbols is
	
	port
	(
		-- Input ports
		index : in integer range 0 to 4;--index : in integer range 0 to 10;
		x_symbol : in integer range 0 to hsymbol;
		y_symbol : in integer range 0 to vsymbol;
		-- Output ports
		rgb_color : out std_logic_vector(2 downto 0) 
	);
end rom_symbols;

architecture lista of rom_symbols is
	
	constant laranja_pou : matrix_symbol :=(
			
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","011","111","111","111","111","111","111","111","110","110","110","111","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","111","111","111","111","111","111","111","111","111","110","110","100","110","111","111","111","111","111","111","111","101","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","111","111","111","111","111","111","111","111","111","110","100","100","100","100","110","111","111","111","111","111","111","111","101","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","100","100","100","100","110","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","011","111","111","111","111","110","110","110","111","111","111","111","100","100","100","100","111","111","111","111","110","110","110","111","111","111","101","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","111","111","111","111","110","110","110","100","110","111","111","111","110","100","100","110","111","111","111","111","100","100","100","110","111","111","111","001","001","001","001","001","001"),
			("001","001","001","001","001","001","011","111","111","111","111","110","100","110","100","100","111","111","111","110","100","110","110","111","111","111","110","100","100","100","110","111","111","111","001","001","001","001","001","001"),
			("001","001","001","001","001","011","111","111","111","111","111","100","110","110","100","100","100","111","111","111","100","100","110","111","111","110","100","100","110","100","100","110","111","111","111","001","001","001","001","001"),
			("001","001","001","001","001","011","111","111","111","111","111","110","100","110","100","100","100","111","111","111","110","100","111","111","111","110","100","100","100","100","110","110","111","111","111","111","001","001","001","001"),
			("001","001","001","001","001","111","111","111","111","111","111","111","110","110","110","100","100","110","111","111","110","110","111","111","110","100","100","100","100","110","110","111","111","111","111","111","001","001","001","001"),
			("001","001","001","001","011","111","111","111","111","111","111","111","111","111","110","110","100","100","110","111","111","110","111","111","100","100","100","110","110","111","111","111","111","111","111","111","001","001","001","001"),
			("001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","110","100","110","110","111","111","111","110","100","110","110","111","111","111","111","111","111","111","111","111","111","001","001","001"),
			("001","001","001","001","111","111","111","111","110","110","110","110","111","111","111","111","111","111","110","110","111","111","111","100","110","111","111","111","111","111","110","110","110","110","111","111","111","001","001","001"),
			("001","001","001","001","111","111","111","110","100","100","100","100","110","110","110","111","111","111","110","111","111","111","111","110","111","111","111","110","110","100","100","100","100","100","110","111","111","001","001","001"),
			("001","001","001","001","111","111","110","110","100","100","100","100","100","100","100","100","110","110","111","111","111","111","111","110","110","110","100","100","100","100","100","100","100","100","110","110","111","001","001","001"),
			("001","001","001","001","111","111","110","110","110","110","110","100","100","100","110","110","111","111","111","111","111","111","111","111","110","110","110","100","100","100","100","100","100","100","110","111","111","001","001","001"),
			("001","001","001","001","111","111","111","110","110","110","110","110","110","111","111","111","111","111","110","110","111","111","111","110","111","111","111","111","111","110","110","100","100","110","111","111","111","001","001","001"),
			("001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","110","100","110","111","111","111","111","110","110","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001"),
			("001","001","001","001","111","111","111","111","111","111","111","111","111","111","110","100","100","100","110","111","110","110","111","110","100","100","110","110","111","111","111","111","111","111","111","111","001","001","001","001"),
			("001","001","001","001","111","111","110","111","111","111","111","111","110","110","100","100","100","110","111","111","110","110","111","111","110","100","100","100","110","111","111","111","111","111","111","111","001","001","001","001"),
			("001","001","001","001","111","111","110","111","111","111","111","110","100","100","100","100","100","111","111","111","110","100","111","111","110","100","110","110","110","110","110","111","111","111","111","111","001","001","001","001"),
			("001","001","001","001","001","111","110","110","111","111","110","100","100","100","100","100","110","111","111","110","100","100","111","111","111","110","110","110","100","100","100","110","111","111","111","111","001","001","001","001"),
			("001","001","001","001","001","111","100","110","110","111","110","100","100","100","100","100","111","111","111","110","100","100","110","111","111","110","110","100","100","100","110","111","111","111","111","111","001","001","001","001"),
			("001","001","001","001","001","001","111","110","110","111","111","110","100","100","100","111","111","111","111","110","110","100","110","111","111","111","110","100","100","100","110","111","111","110","110","001","001","001","001","001"),
			("001","001","001","001","001","001","111","101","110","110","111","110","110","100","110","111","111","111","111","110","110","110","110","111","111","111","111","100","100","110","110","111","110","110","111","001","001","001","001","001"),
			("001","001","001","001","001","001","001","101","100","110","110","111","111","111","111","111","111","111","111","100","100","110","110","110","111","111","111","111","110","110","111","111","110","100","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","101","100","110","110","111","111","111","111","111","111","111","100","100","110","100","110","111","111","111","111","111","111","110","110","100","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","011","001","100","110","110","111","111","111","111","111","111","100","100","110","100","111","111","111","111","111","111","110","110","100","011","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","011","100","100","100","110","110","111","111","111","111","111","110","110","111","111","111","111","111","110","110","100","100","000","011","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","100","100","110","110","110","110","111","111","111","111","111","111","111","110","100","100","100","100","001","011","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","011","100","100","100","100","110","110","110","110","110","110","110","100","100","100","100","101","001","011","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","011","001","100","100","100","100","100","100","100","100","100","100","100","100","001","011","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001")
	);





	
	
	
		constant maca_pou : matrix_symbol :=(
		
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","010","011","010","000","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","010","010","010","000","000","000","010","010","010","011","011","011","011","010","010","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","000","011","111","111","111","111","111","111","111","111","011","010","010","010","010","010","010","010","010","010","011","010","010","010","000","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","000","011","111","111","111","110","110","110","110","111","111","111","110","010","010","010","010","010","010","010","010","010","010","010","010","010","000","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","011","111","111","010","010","110","110","110","110","110","111","110","110","010","010","010","010","010","010","010","010","010","010","010","010","010","010","001","001","001","001","001","001"),
			("001","001","001","001","001","001","011","111","111","010","010","110","111","111","111","111","111","111","111","110","110","010","010","010","010","010","010","010","010","010","010","010","010","010","000","001","001","001","001","001"),
			("001","001","001","001","000","011","111","011","111","111","111","111","111","111","111","111","111","111","111","111","110","110","010","010","010","010","010","010","010","010","010","010","010","010","000","000","001","001","001","001"),
			("001","001","001","001","000","011","011","010","010","111","111","111","111","111","111","111","111","111","111","111","111","110","110","010","010","010","010","010","010","010","010","010","010","010","010","000","001","001","001","001"),
			("001","001","001","001","011","011","010","010","010","111","111","110","111","111","111","111","111","111","110","110","110","110","110","110","010","010","010","010","010","010","010","010","010","010","010","000","001","001","001","001"),
			("001","001","001","011","011","011","010","110","110","111","111","110","111","111","111","111","111","111","110","110","110","110","110","110","010","010","010","010","010","010","010","010","010","010","010","010","001","001","001","001"),
			("001","001","001","011","011","011","110","110","110","110","110","110","110","110","111","111","111","110","110","110","110","110","110","110","010","010","010","010","010","010","010","010","010","010","010","010","001","001","001","001"),
			("001","001","001","001","010","011","010","010","110","110","111","111","110","110","110","110","110","110","110","110","110","110","110","010","010","010","010","010","010","010","010","010","010","010","010","010","000","001","001","001"),
			("001","001","001","011","011","010","010","010","110","110","111","111","110","110","110","110","110","110","110","110","110","110","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","001","001","001"),
			("001","001","001","011","011","010","010","010","110","110","111","110","110","110","110","110","110","110","110","110","110","110","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","001","001","001"),
			("001","001","001","011","011","010","010","110","010","110","110","110","110","110","110","110","110","110","110","110","110","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","001","001","001"),
			("001","001","001","001","010","010","010","110","010","010","110","110","110","110","110","110","110","110","110","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","011","001","001","001","001"),
			("001","001","001","001","010","010","010","010","010","010","010","010","110","110","110","110","010","110","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","011","001","001","001","001"),
			("001","001","001","011","010","011","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","011","001","001","001","001"),
			("001","001","001","011","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","011","001","001","001","001"),
			("001","001","001","011","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","011","001","001","001","001"),
			("001","001","001","011","011","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","011","011","001","001","001","001"),
			("001","001","001","001","011","010","011","011","011","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","011","011","001","001","001","001","001"),
			("001","001","001","001","001","000","010","011","011","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","011","011","001","001","001","001","001"),
			("001","001","001","001","001","001","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","011","011","011","001","001","001","001","001"),
			("001","001","001","001","001","001","001","010","010","010","010","011","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","011","011","011","001","001","001","001","001"),
			("001","001","001","001","001","001","001","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","111","011","011","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","011","011","011","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","011","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","111","011","011","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","011","111","011","010","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","011","011","011","010","010","010","010","010","010","010","010","010","010","010","010","011","011","111","011","011","011","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","011","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","011","011","011","011","010","011","011","011","011","010","010","010","010","011","011","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001")
	);




	
	
	constant pera_pou : matrix_symbol :=(
			
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","101","111","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","111","111","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","011","011","010","000","000","000","111","111","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","011","000","010","110","111","111","011","111","111","111","111","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","010","110","110","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","010","010","110","110","110","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","010","010","110","110","111","111","111","111","111","111","111","011","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","010","010","110","110","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","011","000","000","000","000","010","010","110","110","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","010","010","110","110","110","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","011","000","000","000","000","000","010","010","010","110","110","110","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","000","000","010","010","000","010","010","010","110","110","110","110","111","111","111","111","111","111","111","111","111","011","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","000","000","010","010","110","010","010","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","011","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","000","000","000","000","010","110","010","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","011","000","000","000","000","000","010","010","010","010","110","110","110","111","111","110","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001"),
			("001","001","001","001","001","001","000","000","000","000","000","000","000","010","010","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","001","001","001","001","001"),
			("001","001","001","001","001","001","000","000","000","000","000","000","000","000","010","010","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001"),
			("001","001","001","001","001","001","000","000","000","000","000","000","000","000","010","010","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001"),
			("001","001","001","001","011","000","000","000","000","000","000","000","000","000","010","010","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001"),
			("001","001","001","001","011","000","000","000","000","000","000","000","000","000","010","010","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001"),
			("001","001","001","001","001","000","000","000","000","000","000","000","000","000","010","010","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001"),
			("001","001","001","001","001","000","000","000","000","000","000","000","000","000","010","010","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001"),
			("001","001","001","001","001","000","000","000","000","000","000","000","000","010","010","010","010","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001"),
			("001","001","001","001","001","000","000","000","000","000","000","000","000","000","010","010","010","010","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","011","001","001","001","001","001"),
			("001","001","001","001","011","000","000","000","000","000","000","000","000","000","010","000","010","010","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001"),
			("001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","010","010","010","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","011","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","010","010","010","110","110","110","110","110","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","010","010","010","010","110","110","110","110","110","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","010","010","110","110","110","110","110","110","111","111","111","111","111","111","111","011","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","010","010","010","110","110","110","110","110","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","010","010","110","110","110","110","110","111","111","111","111","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","010","010","010","110","111","111","111","011","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001")
	);






	
	
	constant bola_pou : matrix_symbol :=(
	
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","011","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","000","000","000","001","000","011","111","111","111","111","111","111","111","001","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","000","000","000","001","001","011","111","111","111","111","111","111","111","111","111","000","001","001","000","000","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","000","000","000","000","001","001","001","111","111","111","111","111","111","111","111","111","111","111","001","001","000","000","000","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","000","000","000","000","001","001","111","111","111","111","111","111","111","111","111","111","111","111","001","000","000","000","000","000","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","011","001","000","000","000","000","000","001","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","000","000","000","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","111","001","000","000","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","001","000","000","000","011","001","001","001","001","001","001"),
			("001","001","001","001","001","111","111","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","000","011","111","001","001","001","001","001"),
			("001","001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","001","001","001","001"),
			("001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001"),
			("001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","011","011","011","011","011","011","011","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001"),
			("001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","000","011","111","011","011","011","000","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001"),
			("001","001","001","011","111","111","111","111","111","111","111","111","111","111","111","111","001","000","011","111","111","111","111","001","001","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001"),
			("001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","001","001","001","001","001","001","000","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001"),
			("001","001","001","111","111","011","111","111","111","111","111","111","111","111","111","111","000","000","000","001","001","001","001","000","000","011","111","111","111","111","111","111","111","111","111","111","111","001","001","001"),
			("001","001","001","111","000","000","111","111","111","111","111","111","111","111","111","001","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","001","111","011","001","001"),
			("001","001","001","001","000","000","011","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","111","111","111","111","111","111","111","111","111","000","001","001","001","001"),
			("001","001","001","000","000","000","000","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","000","000","011","111","111","111","111","111","111","111","001","000","000","001","001","001"),
			("001","001","001","000","000","000","000","000","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","000","000","001","111","111","111","111","111","111","111","011","000","000","000","001","001","001"),
			("001","001","001","000","000","000","000","000","001","111","111","111","111","111","111","111","111","000","000","000","000","000","000","000","011","111","111","111","111","111","111","111","011","000","000","000","000","001","001","001"),
			("001","001","001","001","000","000","000","000","000","111","111","111","111","111","111","111","111","111","001","000","000","000","000","111","111","111","111","111","111","111","111","111","001","000","000","000","000","001","001","001"),
			("001","001","001","001","000","000","000","000","001","111","111","111","111","111","111","111","111","111","111","001","000","001","111","111","111","111","111","111","111","111","111","111","001","000","000","000","000","001","001","001"),
			("001","001","001","001","000","000","000","000","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","000","000","000","001","001","001","001"),
			("001","001","001","001","001","000","000","000","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","000","000","000","001","001","001","001"),
			("001","001","001","001","001","000","000","000","001","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","000","000","001","001","001","001","001"),
			("001","001","001","001","001","001","001","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","001","001","001","001","001"),
			("001","001","001","001","001","001","001","011","011","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","011","111","111","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","111","111","011","011","111","111","111","111","111","111","111","011","011","111","111","111","111","111","111","111","011","111","111","011","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","011","111","011","011","111","111","011","011","001","000","000","000","001","011","011","111","111","111","011","111","111","011","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","011","111","111","001","000","000","000","000","000","000","000","000","000","000","001","011","111","111","111","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","111","001","000","000","000","000","000","000","000","000","000","000","000","011","111","011","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","011","001","000","000","000","000","000","000","000","000","000","001","011","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001")
	);




	
	constant bomba_pou : matrix_symbol :=(
	
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","111","111","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","001","001","001","001","000","000","001","001","001","001","001","001","001","110","110","101","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","011","111","111","111","111","111","111","011","001","000","000","000","001","001","001","001","001","001","001","111","111","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","011","111","111","111","111","111","111","111","111","111","011","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","111","111","111","111","111","111","111","111","111","111","111","111","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","000","000","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","111","011","000","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","000","011","111","011","011","111","111","111","111","111","111","111","111","111","111","111","111","111","111","000","000","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","000","000","011","011","011","011","011","011","011","011","011","111","111","111","111","111","111","111","111","111","011","000","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","000","000","000","001","001","011","011","011","011","011","011","011","011","011","011","011","011","111","111","111","111","011","000","000","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","000","001","001","011","011","001","001","001","001","001","011","011","011","011","011","011","011","011","111","111","111","001","000","000","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","000","011","011","111","011","001","001","001","001","001","001","001","001","001","001","011","011","011","011","011","011","000","000","000","000","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","000","001","001","011","001","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001","011","001","000","000","000","000","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","000","001","001","001","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","000","000","001","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","000","000","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","000","001","001","000","000","000","000","000","000","000","000","000","000","000","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001"),
			("001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001","001")
	);




											
begin

	rgb_color <= laranja_pou(y_symbol,x_symbol) 				when index = 0 else
					  maca_pou(y_symbol,x_symbol) 					when index = 1 else
					  pera_pou(y_symbol,x_symbol) 					when index = 2 else
					  bola_pou(y_symbol,x_symbol) 					when index = 3 else
					  bomba_pou(y_symbol,x_symbol) 					when index = 4 else
					  "000";
end lista;
library ieee;
use ieee.std_logic_1164.all;
library work;
use work.vga_package.all;

entity rom_num is
	
	port
	(
		-- Input ports
		index : in integer range 0 to 9;
		x_num : in integer range 0 to hnum;
		y_num : in integer range 0 to vnum;
		-- Output ports
		rgb_num : out std_logic_vector(2 downto 0) 
	);
end rom_num;

architecture lista of rom_num is
	
	constant zero : matrix_num :=(
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","000","000","000","000","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","000","000","000","000","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","000","000","000","000","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","000","000","000","000","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","000","000","000","000","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","000","000","000","000","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010")
	);





	
	constant um : matrix_num :=(
	
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010")
	);




	constant dois : matrix_num :=(
	
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010")
	);



	constant tres : matrix_num :=(
	
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010")
	);



	constant quatro : matrix_num :=(
	
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010")
	);



	constant cinco : matrix_num :=(
	
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010")
	);



	constant seis : matrix_num :=(
		
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010")
	);



	constant sete : matrix_num :=(
	
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010")
	);



	constant oito : matrix_num :=(
	
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010")
	);







	constant nove : matrix_num :=(
	
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010","010","010","010","010","010","010","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010"),
			("010","010","010","010","010","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","000","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010"),
			("010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010","010")
	);









											
begin

	rgb_num <= zero(y_num,x_num) 				when index = 0 else
					  um(y_num,x_num) 				when index = 1 else
					  dois(y_num,x_num) 				when index = 2 else
					  tres(y_num,x_num) 				when index = 3 else
					  quatro(y_num,x_num) 			when index = 4 else
					  cinco(y_num,x_num) 			when index = 5 else
					  seis(y_num,x_num) 				when index = 6 else
					  sete(y_num,x_num) 				when index = 7 else
					  oito(y_num,x_num) 				when index = 8 else
					  nove(y_num,x_num) 				when index = 9 else
						"000";
end lista;